`ifndef MEM_SV
`define MEM_SV

module mem(input  logic        i_clk,
           input  logic        i_reset,
           input  logic [9:0 ] address,
           output logic [31:0] o_data
           );

logic [31:0] mem [0:1023] = '{// T_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F
                              32'hc66363a5, 32'hf87c7c84, 32'hee777799, 32'hf67b7b8d, 32'hfff2f20d, 32'hd66b6bbd, 32'hde6f6fb1, 32'h91c5c554, 32'h60303050, 32'h02010103, 32'hce6767a9, 32'h562b2b7d, 32'he7fefe19, 32'hb5d7d762, 32'h4dababe6, 32'hec76769a,
                              32'h8fcaca45, 32'h1f82829d, 32'h89c9c940, 32'hfa7d7d87, 32'heffafa15, 32'hb25959eb, 32'h8e4747c9, 32'hfbf0f00b, 32'h41adadec, 32'hb3d4d467, 32'h5fa2a2fd, 32'h45afafea, 32'h239c9cbf, 32'h53a4a4f7, 32'he4727296, 32'h9bc0c05b,
                              32'h75b7b7c2, 32'he1fdfd1c, 32'h3d9393ae, 32'h4c26266a, 32'h6c36365a, 32'h7e3f3f41, 32'hf5f7f702, 32'h83cccc4f, 32'h6834345c, 32'h51a5a5f4, 32'hd1e5e534, 32'hf9f1f108, 32'he2717193, 32'habd8d873, 32'h62313153, 32'h2a15153f,
                              32'h0804040c, 32'h95c7c752, 32'h46232365, 32'h9dc3c35e, 32'h30181828, 32'h379696a1, 32'h0a05050f, 32'h2f9a9ab5, 32'h0e070709, 32'h24121236, 32'h1b80809b, 32'hdfe2e23d, 32'hcdebeb26, 32'h4e272769, 32'h7fb2b2cd, 32'hea75759f,
                              32'h1209091b, 32'h1d83839e, 32'h582c2c74, 32'h341a1a2e, 32'h361b1b2d, 32'hdc6e6eb2, 32'hb45a5aee, 32'h5ba0a0fb, 32'ha45252f6, 32'h763b3b4d, 32'hb7d6d661, 32'h7db3b3ce, 32'h5229297b, 32'hdde3e33e, 32'h5e2f2f71, 32'h13848497,
                              32'ha65353f5, 32'hb9d1d168, 32'h00000000, 32'hc1eded2c, 32'h40202060, 32'he3fcfc1f, 32'h79b1b1c8, 32'hb65b5bed, 32'hd46a6abe, 32'h8dcbcb46, 32'h67bebed9, 32'h7239394b, 32'h944a4ade, 32'h984c4cd4, 32'hb05858e8, 32'h85cfcf4a,
                              32'hbbd0d06b, 32'hc5efef2a, 32'h4faaaae5, 32'hedfbfb16, 32'h864343c5, 32'h9a4d4dd7, 32'h66333355, 32'h11858594, 32'h8a4545cf, 32'he9f9f910, 32'h04020206, 32'hfe7f7f81, 32'ha05050f0, 32'h783c3c44, 32'h259f9fba, 32'h4ba8a8e3,
                              32'ha25151f3, 32'h5da3a3fe, 32'h804040c0, 32'h058f8f8a, 32'h3f9292ad, 32'h219d9dbc, 32'h70383848, 32'hf1f5f504, 32'h63bcbcdf, 32'h77b6b6c1, 32'hafdada75, 32'h42212163, 32'h20101030, 32'he5ffff1a, 32'hfdf3f30e, 32'hbfd2d26d,
                              32'h81cdcd4c, 32'h180c0c14, 32'h26131335, 32'hc3ecec2f, 32'hbe5f5fe1, 32'h359797a2, 32'h884444cc, 32'h2e171739, 32'h93c4c457, 32'h55a7a7f2, 32'hfc7e7e82, 32'h7a3d3d47, 32'hc86464ac, 32'hba5d5de7, 32'h3219192b, 32'he6737395,
                              32'hc06060a0, 32'h19818198, 32'h9e4f4fd1, 32'ha3dcdc7f, 32'h44222266, 32'h542a2a7e, 32'h3b9090ab, 32'h0b888883, 32'h8c4646ca, 32'hc7eeee29, 32'h6bb8b8d3, 32'h2814143c, 32'ha7dede79, 32'hbc5e5ee2, 32'h160b0b1d, 32'haddbdb76,
                              32'hdbe0e03b, 32'h64323256, 32'h743a3a4e, 32'h140a0a1e, 32'h924949db, 32'h0c06060a, 32'h4824246c, 32'hb85c5ce4, 32'h9fc2c25d, 32'hbdd3d36e, 32'h43acacef, 32'hc46262a6, 32'h399191a8, 32'h319595a4, 32'hd3e4e437, 32'hf279798b,
                              32'hd5e7e732, 32'h8bc8c843, 32'h6e373759, 32'hda6d6db7, 32'h018d8d8c, 32'hb1d5d564, 32'h9c4e4ed2, 32'h49a9a9e0, 32'hd86c6cb4, 32'hac5656fa, 32'hf3f4f407, 32'hcfeaea25, 32'hca6565af, 32'hf47a7a8e, 32'h47aeaee9, 32'h10080818,
                              32'h6fbabad5, 32'hf0787888, 32'h4a25256f, 32'h5c2e2e72, 32'h381c1c24, 32'h57a6a6f1, 32'h73b4b4c7, 32'h97c6c651, 32'hcbe8e823, 32'ha1dddd7c, 32'he874749c, 32'h3e1f1f21, 32'h964b4bdd, 32'h61bdbddc, 32'h0d8b8b86, 32'h0f8a8a85,
                              32'he0707090, 32'h7c3e3e42, 32'h71b5b5c4, 32'hcc6666aa, 32'h904848d8, 32'h06030305, 32'hf7f6f601, 32'h1c0e0e12, 32'hc26161a3, 32'h6a35355f, 32'hae5757f9, 32'h69b9b9d0, 32'h17868691, 32'h99c1c158, 32'h3a1d1d27, 32'h279e9eb9,
                              32'hd9e1e138, 32'hebf8f813, 32'h2b9898b3, 32'h22111133, 32'hd26969bb, 32'ha9d9d970, 32'h078e8e89, 32'h339494a7, 32'h2d9b9bb6, 32'h3c1e1e22, 32'h15878792, 32'hc9e9e920, 32'h87cece49, 32'haa5555ff, 32'h50282878, 32'ha5dfdf7a,
                              32'h038c8c8f, 32'h59a1a1f8, 32'h09898980, 32'h1a0d0d17, 32'h65bfbfda, 32'hd7e6e631, 32'h844242c6, 32'hd06868b8, 32'h824141c3, 32'h299999b0, 32'h5a2d2d77, 32'h1e0f0f11, 32'h7bb0b0cb, 32'ha85454fc, 32'h6dbbbbd6, 32'h2c16163a,
                              // S_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F                              
										32'h63000000, 32'h7c000000, 32'h77000000, 32'h7b000000, 32'hf2000000, 32'h6b000000, 32'h6f000000, 32'hc5000000, 32'h30000000, 32'h01000000, 32'h67000000, 32'h2b000000, 32'hfe000000, 32'hd7000000, 32'hab000000, 32'h76000000, 
                              32'hca000000, 32'h82000000, 32'hc9000000, 32'h7d000000, 32'hfa000000, 32'h59000000, 32'h47000000, 32'hf0000000, 32'had000000, 32'hd4000000, 32'ha2000000, 32'haf000000, 32'h9c000000, 32'ha4000000, 32'h72000000, 32'hc0000000, 
                              32'hb7000000, 32'hfd000000, 32'h93000000, 32'h26000000, 32'h36000000, 32'h3f000000, 32'hf7000000, 32'hcc000000, 32'h34000000, 32'ha5000000, 32'he5000000, 32'hf1000000, 32'h71000000, 32'hd8000000, 32'h31000000, 32'h15000000, 
                              32'h04000000, 32'hc7000000, 32'h23000000, 32'hc3000000, 32'h18000000, 32'h96000000, 32'h05000000, 32'h9a000000, 32'h07000000, 32'h12000000, 32'h80000000, 32'he2000000, 32'heb000000, 32'h27000000, 32'hb2000000, 32'h75000000, 
                              32'h09000000, 32'h83000000, 32'h2c000000, 32'h1a000000, 32'h1b000000, 32'h6e000000, 32'h5a000000, 32'ha0000000, 32'h52000000, 32'h3b000000, 32'hd6000000, 32'hb3000000, 32'h29000000, 32'he3000000, 32'h2f000000, 32'h84000000, 
                              32'h53000000, 32'hd1000000, 32'h00000000, 32'hed000000, 32'h20000000, 32'hfc000000, 32'hb1000000, 32'h5b000000, 32'h6a000000, 32'hcb000000, 32'hbe000000, 32'h39000000, 32'h4a000000, 32'h4c000000, 32'h58000000, 32'hcf000000, 
                              32'hd0000000, 32'hef000000, 32'haa000000, 32'hfb000000, 32'h43000000, 32'h4d000000, 32'h33000000, 32'h85000000, 32'h45000000, 32'hf9000000, 32'h02000000, 32'h7f000000, 32'h50000000, 32'h3c000000, 32'h9f000000, 32'ha8000000, 
                              32'h51000000, 32'ha3000000, 32'h40000000, 32'h8f000000, 32'h92000000, 32'h9d000000, 32'h38000000, 32'hf5000000, 32'hbc000000, 32'hb6000000, 32'hda000000, 32'h21000000, 32'h10000000, 32'hff000000, 32'hf3000000, 32'hd2000000, 
                              32'hcd000000, 32'h0c000000, 32'h13000000, 32'hec000000, 32'h5f000000, 32'h97000000, 32'h44000000, 32'h17000000, 32'hc4000000, 32'ha7000000, 32'h7e000000, 32'h3d000000, 32'h64000000, 32'h5d000000, 32'h19000000, 32'h73000000, 
                              32'h60000000, 32'h81000000, 32'h4f000000, 32'hdc000000, 32'h22000000, 32'h2a000000, 32'h90000000, 32'h88000000, 32'h46000000, 32'hee000000, 32'hb8000000, 32'h14000000, 32'hde000000, 32'h5e000000, 32'h0b000000, 32'hdb000000, 
                              32'he0000000, 32'h32000000, 32'h3a000000, 32'h0a000000, 32'h49000000, 32'h06000000, 32'h24000000, 32'h5c000000, 32'hc2000000, 32'hd3000000, 32'hac000000, 32'h62000000, 32'h91000000, 32'h95000000, 32'he4000000, 32'h79000000, 
                              32'he7000000, 32'hc8000000, 32'h37000000, 32'h6d000000, 32'h8d000000, 32'hd5000000, 32'h4e000000, 32'ha9000000, 32'h6c000000, 32'h56000000, 32'hf4000000, 32'hea000000, 32'h65000000, 32'h7a000000, 32'hae000000, 32'h08000000, 
                              32'hba000000, 32'h78000000, 32'h25000000, 32'h2e000000, 32'h1c000000, 32'ha6000000, 32'hb4000000, 32'hc6000000, 32'he8000000, 32'hdd000000, 32'h74000000, 32'h1f000000, 32'h4b000000, 32'hbd000000, 32'h8b000000, 32'h8a000000, 
                              32'h70000000, 32'h3e000000, 32'hb5000000, 32'h66000000, 32'h48000000, 32'h03000000, 32'hf6000000, 32'h0e000000, 32'h61000000, 32'h35000000, 32'h57000000, 32'hb9000000, 32'h86000000, 32'hc1000000, 32'h1d000000, 32'h9e000000, 
                              32'he1000000, 32'hf8000000, 32'h98000000, 32'h11000000, 32'h69000000, 32'hd9000000, 32'h8e000000, 32'h94000000, 32'h9b000000, 32'h1e000000, 32'h87000000, 32'he9000000, 32'hce000000, 32'h55000000, 32'h28000000, 32'hdf000000, 
                              32'h8c000000, 32'ha1000000, 32'h89000000, 32'h0d000000, 32'hbf000000, 32'he6000000, 32'h42000000, 32'h68000000, 32'h41000000, 32'h99000000, 32'h2d000000, 32'h0f000000, 32'hb0000000, 32'h54000000, 32'hbb000000, 32'h16000000,
                              // Inv_T_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F                              
							32'h51f4a750, 32'h7e416553, 32'h1a17a4c3, 32'h3a275e96, 32'h3bab6bcb, 32'h1f9d45f1, 32'hacfa58ab, 32'h4be30393, 32'h2030fa55, 32'had766df6, 32'h88cc7691, 32'hf5024c25, 32'h4fe5d7fc, 32'hc52acbd7, 32'h26354480, 32'hb562a38f,
                              32'hdeb15a49, 32'h25ba1b67, 32'h45ea0e98, 32'h5dfec0e1, 32'hc32f7502, 32'h814cf012, 32'h8d4697a3, 32'h6bd3f9c6, 32'h038f5fe7, 32'h15929c95, 32'hbf6d7aeb, 32'h955259da, 32'hd4be832d, 32'h587421d3, 32'h49e06929, 32'h8ec9c844,
                              32'h75c2896a, 32'hf48e7978, 32'h99583e6b, 32'h27b971dd, 32'hbee14fb6, 32'hf088ad17, 32'hc920ac66, 32'h7dce3ab4, 32'h63df4a18, 32'he51a3182, 32'h97513360, 32'h62537f45, 32'hb16477e0, 32'hbb6bae84, 32'hfe81a01c, 32'hf9082b94,
                              32'h70486858, 32'h8f45fd19, 32'h94de6c87, 32'h527bf8b7, 32'hab73d323, 32'h724b02e2, 32'he31f8f57, 32'h6655ab2a, 32'hb2eb2807, 32'h2fb5c203, 32'h86c57b9a, 32'hd33708a5, 32'h302887f2, 32'h23bfa5b2, 32'h02036aba, 32'hed16825c,
                              32'h8acf1c2b, 32'ha779b492, 32'hf307f2f0, 32'h4e69e2a1, 32'h65daf4cd, 32'h0605bed5, 32'hd134621f, 32'hc4a6fe8a, 32'h342e539d, 32'ha2f355a0, 32'h058ae132, 32'ha4f6eb75, 32'h0b83ec39, 32'h4060efaa, 32'h5e719f06, 32'hbd6e1051,
                              32'h3e218af9, 32'h96dd063d, 32'hdd3e05ae, 32'h4de6bd46, 32'h91548db5, 32'h71c45d05, 32'h0406d46f, 32'h605015ff, 32'h1998fb24, 32'hd6bde997, 32'h894043cc, 32'h67d99e77, 32'hb0e842bd, 32'h07898b88, 32'he7195b38, 32'h79c8eedb,
                              32'ha17c0a47, 32'h7c420fe9, 32'hf8841ec9, 32'h00000000, 32'h09808683, 32'h322bed48, 32'h1e1170ac, 32'h6c5a724e, 32'hfd0efffb, 32'h0f853856, 32'h3daed51e, 32'h362d3927, 32'h0a0fd964, 32'h685ca621, 32'h9b5b54d1, 32'h24362e3a,
                              32'h0c0a67b1, 32'h9357e70f, 32'hb4ee96d2, 32'h1b9b919e, 32'h80c0c54f, 32'h61dc20a2, 32'h5a774b69, 32'h1c121a16, 32'he293ba0a, 32'hc0a02ae5, 32'h3c22e043, 32'h121b171d, 32'h0e090d0b, 32'hf28bc7ad, 32'h2db6a8b9, 32'h141ea9c8,
                              32'h57f11985, 32'haf75074c, 32'hee99ddbb, 32'ha37f60fd, 32'hf701269f, 32'h5c72f5bc, 32'h44663bc5, 32'h5bfb7e34, 32'h8b432976, 32'hcb23c6dc, 32'hb6edfc68, 32'hb8e4f163, 32'hd731dcca, 32'h42638510, 32'h13972240, 32'h84c61120,
                              32'h854a247d, 32'hd2bb3df8, 32'haef93211, 32'hc729a16d, 32'h1d9e2f4b, 32'hdcb230f3, 32'h0d8652ec, 32'h77c1e3d0, 32'h2bb3166c, 32'ha970b999, 32'h119448fa, 32'h47e96422, 32'ha8fc8cc4, 32'ha0f03f1a, 32'h567d2cd8, 32'h223390ef,
                              32'h87494ec7, 32'hd938d1c1, 32'h8ccaa2fe, 32'h98d40b36, 32'ha6f581cf, 32'ha57ade28, 32'hdab78e26, 32'h3fadbfa4, 32'h2c3a9de4, 32'h5078920d, 32'h6a5fcc9b, 32'h547e4662, 32'hf68d13c2, 32'h90d8b8e8, 32'h2e39f75e, 32'h82c3aff5,
                              32'h9f5d80be, 32'h69d0937c, 32'h6fd52da9, 32'hcf2512b3, 32'hc8ac993b, 32'h10187da7, 32'he89c636e, 32'hdb3bbb7b, 32'hcd267809, 32'h6e5918f4, 32'hec9ab701, 32'h834f9aa8, 32'he6956e65, 32'haaffe67e, 32'h21bccf08, 32'hef15e8e6,
                              32'hbae79bd9, 32'h4a6f36ce, 32'hea9f09d4, 32'h29b07cd6, 32'h31a4b2af, 32'h2a3f2331, 32'hc6a59430, 32'h35a266c0, 32'h744ebc37, 32'hfc82caa6, 32'he090d0b0, 32'h33a7d815, 32'hf104984a, 32'h41ecdaf7, 32'h7fcd500e, 32'h1791f62f,
                              32'h764dd68d, 32'h43efb04d, 32'hccaa4d54, 32'he49604df, 32'h9ed1b5e3, 32'h4c6a881b, 32'hc12c1fb8, 32'h4665517f, 32'h9d5eea04, 32'h018c355d, 32'hfa877473, 32'hfb0b412e, 32'hb3671d5a, 32'h92dbd252, 32'he9105633, 32'h6dd64713,
                              32'h9ad7618c, 32'h37a10c7a, 32'h59f8148e, 32'heb133c89, 32'hcea927ee, 32'hb761c935, 32'he11ce5ed, 32'h7a47b13c, 32'h9cd2df59, 32'h55f2733f, 32'h1814ce79, 32'h73c737bf, 32'h53f7cdea, 32'h5ffdaa5b, 32'hdf3d6f14, 32'h7844db86,
                              32'hcaaff381, 32'hb968c43e, 32'h3824342c, 32'hc2a3405f, 32'h161dc372, 32'hbce2250c, 32'h283c498b, 32'hff0d9541, 32'h39a80171, 32'h080cb3de, 32'hd8b4e49c, 32'h6456c190, 32'h7bcb8461, 32'hd532b670, 32'h486c5c74, 32'hd0b85742,
                              // Inv_S_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E                                                                  
					32'h52000000, 32'h09000000, 32'h6a000000, 32'hd5000000, 32'h30000000, 32'h36000000, 32'ha5000000, 32'h38000000, 32'hbf000000, 32'h40000000, 32'ha3000000, 32'h9e000000, 32'h81000000, 32'hf3000000, 32'hd7000000, 32'hfb000000, 
                              32'h7c000000, 32'he3000000, 32'h39000000, 32'h82000000, 32'h9b000000, 32'h2f000000, 32'hff000000, 32'h87000000, 32'h34000000, 32'h8e000000, 32'h43000000, 32'h44000000, 32'hc4000000, 32'hde000000, 32'he9000000, 32'hcb000000, 
                              32'h54000000, 32'h7b000000, 32'h94000000, 32'h32000000, 32'ha6000000, 32'hc2000000, 32'h23000000, 32'h3d000000, 32'hee000000, 32'h4c000000, 32'h95000000, 32'h0b000000, 32'h42000000, 32'hfa000000, 32'hc3000000, 32'h4e000000, 
                              32'h08000000, 32'h2e000000, 32'ha1000000, 32'h66000000, 32'h28000000, 32'hd9000000, 32'h24000000, 32'hb2000000, 32'h76000000, 32'h5b000000, 32'ha2000000, 32'h49000000, 32'h6d000000, 32'h8b000000, 32'hd1000000, 32'h25000000, 
                              32'h72000000, 32'hf8000000, 32'hf6000000, 32'h64000000, 32'h86000000, 32'h68000000, 32'h98000000, 32'h16000000, 32'hd4000000, 32'ha4000000, 32'h5c000000, 32'hcc000000, 32'h5d000000, 32'h65000000, 32'hb6000000, 32'h92000000, 
                              32'h6c000000, 32'h70000000, 32'h48000000, 32'h50000000, 32'hfd000000, 32'hed000000, 32'hb9000000, 32'hda000000, 32'h5e000000, 32'h15000000, 32'h46000000, 32'h57000000, 32'ha7000000, 32'h8d000000, 32'h9d000000, 32'h84000000, 
                              32'h90000000, 32'hd8000000, 32'hab000000, 32'h00000000, 32'h8c000000, 32'hbc000000, 32'hd3000000, 32'h0a000000, 32'hf7000000, 32'he4000000, 32'h58000000, 32'h05000000, 32'hb8000000, 32'hb3000000, 32'h45000000, 32'h06000000, 
                              32'hd0000000, 32'h2c000000, 32'h1e000000, 32'h8f000000, 32'hca000000, 32'h3f000000, 32'h0f000000, 32'h02000000, 32'hc1000000, 32'haf000000, 32'hbd000000, 32'h03000000, 32'h01000000, 32'h13000000, 32'h8a000000, 32'h6b000000, 
                              32'h3a000000, 32'h91000000, 32'h11000000, 32'h41000000, 32'h4f000000, 32'h67000000, 32'hdc000000, 32'hea000000, 32'h97000000, 32'hf2000000, 32'hcf000000, 32'hce000000, 32'hf0000000, 32'hb4000000, 32'he6000000, 32'h73000000, 
                              32'h96000000, 32'hac000000, 32'h74000000, 32'h22000000, 32'he7000000, 32'had000000, 32'h35000000, 32'h85000000, 32'he2000000, 32'hf9000000, 32'h37000000, 32'he8000000, 32'h1c000000, 32'h75000000, 32'hdf000000, 32'h6e000000, 
                              32'h47000000, 32'hf1000000, 32'h1a000000, 32'h71000000, 32'h1d000000, 32'h29000000, 32'hc5000000, 32'h89000000, 32'h6f000000, 32'hb7000000, 32'h62000000, 32'h0e000000, 32'haa000000, 32'h18000000, 32'hbe000000, 32'h1b000000, 
                              32'hfc000000, 32'h56000000, 32'h3e000000, 32'h4b000000, 32'hc6000000, 32'hd2000000, 32'h79000000, 32'h20000000, 32'h9a000000, 32'hdb000000, 32'hc0000000, 32'hfe000000, 32'h78000000, 32'hcd000000, 32'h5a000000, 32'hf4000000, 
                              32'h1f000000, 32'hdd000000, 32'ha8000000, 32'h33000000, 32'h88000000, 32'h07000000, 32'hc7000000, 32'h31000000, 32'hb1000000, 32'h12000000, 32'h10000000, 32'h59000000, 32'h27000000, 32'h80000000, 32'hec000000, 32'h5f000000, 
                              32'h60000000, 32'h51000000, 32'h7f000000, 32'ha9000000, 32'h19000000, 32'hb5000000, 32'h4a000000, 32'h0d000000, 32'h2d000000, 32'he5000000, 32'h7a000000, 32'h9f000000, 32'h93000000, 32'hc9000000, 32'h9c000000, 32'hef000000, 
                              32'ha0000000, 32'he0000000, 32'h3b000000, 32'h4d000000, 32'hae000000, 32'h2a000000, 32'hf5000000, 32'hb0000000, 32'hc8000000, 32'heb000000, 32'hbb000000, 32'h3c000000, 32'h83000000, 32'h53000000, 32'h99000000, 32'h61000000, 
                              32'h17000000, 32'h2b000000, 32'h04000000, 32'h7e000000, 32'hba000000, 32'h77000000, 32'hd6000000, 32'h26000000, 32'he1000000, 32'h69000000, 32'h14000000, 32'h63000000, 32'h55000000, 32'h21000000, 32'h0c000000, 32'h7d000000
                              };
									
always_comb begin
      if(!i_reset) begin
            o_data = 32'h0;
      end
      else
      begin
            o_data = mem[address];
      end
end		 

endmodule 

`endif