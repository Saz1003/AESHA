`ifndef RC_SV
`define RC_SV

module rc (input [4:0] t, output logic [63:0] rct);

	always_comb begin
		case (t)
			5'b00000: rct = 64'h0000000000000001;
			5'b00001: rct = 64'h0000000000008082;
			5'b00010: rct = 64'h800000000000808A;
			5'b00011: rct = 64'h8000000080008000;
			5'b00100: rct = 64'h000000000000808B;
			5'b00101: rct = 64'h0000000080000001;
			5'b00110: rct = 64'h8000000080008081;
			5'b00111: rct = 64'h8000000000008009;
			5'b01000: rct = 64'h000000000000008A;
			5'b01001: rct = 64'h0000000000000088;
			5'b01010: rct = 64'h0000000080008009;
			5'b01011: rct = 64'h000000008000000A;
			5'b01100: rct = 64'h000000008000808B;
			5'b01101: rct = 64'h800000000000008B;
			5'b01110: rct = 64'h8000000000008089;
			5'b01111: rct = 64'h8000000000008003;
			5'b10000: rct = 64'h8000000000008002;
			5'b10001: rct = 64'h8000000000000080;
			5'b10010: rct = 64'h000000000000800A;
			5'b10011: rct = 64'h800000008000000A;
			5'b10100: rct = 64'h8000000080008081;
			5'b10101: rct = 64'h8000000000008080;
			5'b10110: rct = 64'h0000000080000001;
			5'b10111: rct = 64'h8000000080008008;
			default: rct = 64'h0;
		endcase
	end

endmodule

`endif // RC_SV