`ifndef MEM_SV
`define MEM_SV

module mem(input  logic        i_clk,
           input  logic        i_reset,
           input  logic [9:0 ] address,
           output logic [31:0] o_data
           );

logic [31:0] mem [0:1023] = '{// T_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F
                              32'hc66363a5, 32'hf87c7c84, 32'hee777799, 32'hf67b7b8d, 32'hfff2f20d, 32'hd66b6bbd, 32'hde6f6fb1, 32'h91c5c554, 32'h60303050, 32'h02010103, 32'hce6767a9, 32'h562b2b7d, 32'he7fefe19, 32'hb5d7d762, 32'h4dababe6, 32'hec76769a, 
                              32'h8fcaca45, 32'h1f82829d, 32'h89c9c940, 32'hfa7d7d87, 32'heffafa15, 32'hb25959eb, 32'h8e4747c9, 32'hfbf0f00b, 32'h41adadec, 32'hb3d4d467, 32'h5fa2a2fd, 32'h45afafea, 32'h239c9cbf, 32'h53a4a4f7, 32'he4727296, 32'h9bc0c05b, 
                              32'h75b7b7c2, 32'he1fdfd1c, 32'h3d9393ae, 32'h4c26266a, 32'h6c36365a, 32'h7e3f3f41, 32'hf5f7f702, 32'h83cccc4f, 32'h6834345c, 32'h51a5a5f4, 32'hd1e5e534, 32'hf9f1f108, 32'he2717193, 32'habd8d873, 32'h62313153, 32'h2a15153f, 
                              32'h0804040c, 32'h95c7c752, 32'h46232365, 32'h9dc3c35e, 32'h30181828, 32'h379696a1, 32'h0a05050f, 32'h2f9a9ab5, 32'h0e070709, 32'h24121236, 32'h1b80809b, 32'hdfe2e23d, 32'hcdebeb26, 32'h4e272769, 32'h7fb2b2cd, 32'hea75759f, 
                              32'h1209091b, 32'h1d83839e, 32'h582c2c74, 32'h341a1a2e, 32'h361b1b2d, 32'hdc6e6eb2, 32'hb45a5aee, 32'h5ba0a0fb, 32'ha45252f6, 32'h763b3b4d, 32'hb7d6d661, 32'h7db3b3ce, 32'h5229297b, 32'hdde3e33e, 32'h5e2f2f71, 32'h13848497, 
                              32'ha65353f5, 32'hb9d1d168, 32'h00000000, 32'hc1eded2c, 32'h40202060, 32'he3fcfc1f, 32'h79b1b1c8, 32'hb65b5bed, 32'hd46a6abe, 32'h8dcbcb46, 32'h67bebed9, 32'h7239394b, 32'h944a4ade, 32'h984c4cd4, 32'hb05858e8, 32'h85cfcf4a, 
                              32'hbbd0d06b, 32'hc5efef2a, 32'h4faaaae5, 32'hedfbfb16, 32'h864343c5, 32'h9a4d4dd7, 32'h66333355, 32'h11858594, 32'h8a4545cf, 32'he9f9f910, 32'h04020206, 32'hfe7f7f81, 32'ha05050f0, 32'h783c3c44, 32'h259f9fba, 32'h4ba8a8e3, 
                              32'ha25151f3, 32'h5da3a3fe, 32'h804040c0, 32'h058f8f8a, 32'h3f9292ad, 32'h219d9dbc, 32'h70383848, 32'hf1f5f504, 32'h63bcbcdf, 32'h77b6b6c1, 32'hafdada75, 32'h42212163, 32'h20101030, 32'he5ffff1a, 32'hfdf3f30e, 32'hbfd2d26d, 
                              32'h81cdcd4c, 32'h180c0c14, 32'h26131335, 32'hc3ecec2f, 32'hbe5f5fe1, 32'h359797a2, 32'h884444cc, 32'h2e171739, 32'h93c4c457, 32'h55a7a7f2, 32'hfc7e7e82, 32'h7a3d3d47, 32'hc86464ac, 32'hba5d5de7, 32'h3219192b, 32'he6737395, 
                              32'hc06060a0, 32'h19818198, 32'h9e4f4fd1, 32'ha3dcdc7f, 32'h44222266, 32'h542a2a7e, 32'h3b9090ab, 32'h0b888883, 32'h8c4646ca, 32'hc7eeee29, 32'h6bb8b8d3, 32'h2814143c, 32'ha7dede79, 32'hbc5e5ee2, 32'h160b0b1d, 32'haddbdb76, 
                              32'hdbe0e03b, 32'h64323256, 32'h743a3a4e, 32'h140a0a1e, 32'h924949db, 32'h0c06060a, 32'h4824246c, 32'hb85c5ce4, 32'h9fc2c25d, 32'hbdd3d36e, 32'h43acacef, 32'hc46262a6, 32'h399191a8, 32'h319595a4, 32'hd3e4e437, 32'hf279798b, 
                              32'hd5e7e732, 32'h8bc8c843, 32'h6e373759, 32'hda6d6db7, 32'h018d8d8c, 32'hb1d5d564, 32'h9c4e4ed2, 32'h49a9a9e0, 32'hd86c6cb4, 32'hac5656fa, 32'hf3f4f407, 32'hcfeaea25, 32'hca6565af, 32'hf47a7a8e, 32'h47aeaee9, 32'h10080818, 
                              32'h6fbabad5, 32'hf0787888, 32'h4a25256f, 32'h5c2e2e72, 32'h381c1c24, 32'h57a6a6f1, 32'h73b4b4c7, 32'h97c6c651, 32'hcbe8e823, 32'ha1dddd7c, 32'he874749c, 32'h3e1f1f21, 32'h964b4bdd, 32'h61bdbddc, 32'h0d8b8b86, 32'h0f8a8a85, 
                              32'he0707090, 32'h7c3e3e42, 32'h71b5b5c4, 32'hcc6666aa, 32'h904848d8, 32'h06030305, 32'hf7f6f601, 32'h1c0e0e12, 32'hc26161a3, 32'h6a35355f, 32'hae5757f9, 32'h69b9b9d0, 32'h17868691, 32'h99c1c158, 32'h3a1d1d27, 32'h279e9eb9, 
                              32'hd9e1e138, 32'hebf8f813, 32'h2b9898b3, 32'h22111133, 32'hd26969bb, 32'ha9d9d970, 32'h078e8e89, 32'h339494a7, 32'h2d9b9bb6, 32'h3c1e1e22, 32'h15878792, 32'hc9e9e920, 32'h87cece49, 32'haa5555ff, 32'h50282878, 32'ha5dfdf7a, 
                              32'h038c8c8f, 32'h59a1a1f8, 32'h09898980, 32'h1a0d0d17, 32'h65bfbfda, 32'hd7e6e631, 32'h844242c6, 32'hd06868b8, 32'h824141c3, 32'h299999b0, 32'h5a2d2d77, 32'h1e0f0f11, 32'h7bb0b0cb, 32'ha85454fc, 32'h6dbbbbd6, 32'h2c16163a, 
                              // S_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F                              
					32'h63000000, 32'h7c000000, 32'h77000000, 32'h7b000000, 32'hf2000000, 32'h6b000000, 32'h6f000000, 32'hc5000000, 32'h30000000, 32'h01000000, 32'h67000000, 32'h2b000000, 32'hfe000000, 32'hd7000000, 32'hab000000, 32'h76000000, 
                              32'hca000000, 32'h82000000, 32'hc9000000, 32'h7d000000, 32'hfa000000, 32'h59000000, 32'h47000000, 32'hf0000000, 32'had000000, 32'hd4000000, 32'ha2000000, 32'haf000000, 32'h9c000000, 32'ha4000000, 32'h72000000, 32'hc0000000, 
                              32'hb7000000, 32'hfd000000, 32'h93000000, 32'h26000000, 32'h36000000, 32'h3f000000, 32'hf7000000, 32'hcc000000, 32'h34000000, 32'ha5000000, 32'he5000000, 32'hf1000000, 32'h71000000, 32'hd8000000, 32'h31000000, 32'h15000000, 
                              32'h04000000, 32'hc7000000, 32'h23000000, 32'hc3000000, 32'h18000000, 32'h96000000, 32'h05000000, 32'h9a000000, 32'h07000000, 32'h12000000, 32'h80000000, 32'he2000000, 32'heb000000, 32'h27000000, 32'hb2000000, 32'h75000000, 
                              32'h09000000, 32'h83000000, 32'h2c000000, 32'h1a000000, 32'h1b000000, 32'h6e000000, 32'h5a000000, 32'ha0000000, 32'h52000000, 32'h3b000000, 32'hd6000000, 32'hb3000000, 32'h29000000, 32'he3000000, 32'h2f000000, 32'h84000000, 
                              32'h53000000, 32'hd1000000, 32'h00000000, 32'hed000000, 32'h20000000, 32'hfc000000, 32'hb1000000, 32'h5b000000, 32'h6a000000, 32'hcb000000, 32'hbe000000, 32'h39000000, 32'h4a000000, 32'h4c000000, 32'h58000000, 32'hcf000000, 
                              32'hd0000000, 32'hef000000, 32'haa000000, 32'hfb000000, 32'h43000000, 32'h4d000000, 32'h33000000, 32'h85000000, 32'h45000000, 32'hf9000000, 32'h02000000, 32'h7f000000, 32'h50000000, 32'h3c000000, 32'h9f000000, 32'ha8000000, 
                              32'h51000000, 32'ha3000000, 32'h40000000, 32'h8f000000, 32'h92000000, 32'h9d000000, 32'h38000000, 32'hf5000000, 32'hbc000000, 32'hb6000000, 32'hda000000, 32'h21000000, 32'h10000000, 32'hff000000, 32'hf3000000, 32'hd2000000, 
                              32'hcd000000, 32'h0c000000, 32'h13000000, 32'hec000000, 32'h5f000000, 32'h97000000, 32'h44000000, 32'h17000000, 32'hc4000000, 32'ha7000000, 32'h7e000000, 32'h3d000000, 32'h64000000, 32'h5d000000, 32'h19000000, 32'h73000000, 
                              32'h60000000, 32'h81000000, 32'h4f000000, 32'hdc000000, 32'h22000000, 32'h2a000000, 32'h90000000, 32'h88000000, 32'h46000000, 32'hee000000, 32'hb8000000, 32'h14000000, 32'hde000000, 32'h5e000000, 32'h0b000000, 32'hdb000000, 
                              32'he0000000, 32'h32000000, 32'h3a000000, 32'h0a000000, 32'h49000000, 32'h06000000, 32'h24000000, 32'h5c000000, 32'hc2000000, 32'hd3000000, 32'hac000000, 32'h62000000, 32'h91000000, 32'h95000000, 32'he4000000, 32'h79000000, 
                              32'he7000000, 32'hc8000000, 32'h37000000, 32'h6d000000, 32'h8d000000, 32'hd5000000, 32'h4e000000, 32'ha9000000, 32'h6c000000, 32'h56000000, 32'hf4000000, 32'hea000000, 32'h65000000, 32'h7a000000, 32'hae000000, 32'h08000000, 
                              32'hba000000, 32'h78000000, 32'h25000000, 32'h2e000000, 32'h1c000000, 32'ha6000000, 32'hb4000000, 32'hc6000000, 32'he8000000, 32'hdd000000, 32'h74000000, 32'h1f000000, 32'h4b000000, 32'hbd000000, 32'h8b000000, 32'h8a000000, 
                              32'h70000000, 32'h3e000000, 32'hb5000000, 32'h66000000, 32'h48000000, 32'h03000000, 32'hf6000000, 32'h0e000000, 32'h61000000, 32'h35000000, 32'h57000000, 32'hb9000000, 32'h86000000, 32'hc1000000, 32'h1d000000, 32'h9e000000, 
                              32'he1000000, 32'hf8000000, 32'h98000000, 32'h11000000, 32'h69000000, 32'hd9000000, 32'h8e000000, 32'h94000000, 32'h9b000000, 32'h1e000000, 32'h87000000, 32'he9000000, 32'hce000000, 32'h55000000, 32'h28000000, 32'hdf000000, 
                              32'h8c000000, 32'ha1000000, 32'h89000000, 32'h0d000000, 32'hbf000000, 32'he6000000, 32'h42000000, 32'h68000000, 32'h41000000, 32'h99000000, 32'h2d000000, 32'h0f000000, 32'hb0000000, 32'h54000000, 32'hbb000000, 32'h16000000,
                              // Inv_T_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E             F                              
					32'h51F4A750, 32'h7E416553, 32'h1A17A4C3, 32'h3A275E96, 32'h3BAB6BCB, 32'h1F9D45F1, 32'hACFA58AB, 32'h4BE30393, 32'h2030FA55, 32'hAD766DF6, 32'h88CC7691, 32'hF5024C25, 32'h4FE5D7FC, 32'hC52ACBD7, 32'h26354480, 32'hB562A38F, 
                              32'hDEB15A49, 32'h25BA1B67, 32'h45EA0E98, 32'h5DFEC0E1, 32'hC32F7502, 32'h814CF012, 32'h8D4697A3, 32'h6BD3F9C6, 32'h038F5FE7, 32'h15929C95, 32'hBF6D7AEB, 32'h955259DA, 32'hD4BE832D, 32'h587421D3, 32'h49E06929, 32'h8EC9C844, 
                              32'h75C2896A, 32'hF48E7978, 32'h99583E6B, 32'h27B971DD, 32'hBEE14FB6, 32'hF088AD17, 32'hC920AC66, 32'h7DCE3AB4, 32'h63DF4A18, 32'hE51A3182, 32'h97513360, 32'h62537F45, 32'hB16477E0, 32'hBB6BAE84, 32'hFE81A01C, 32'hF9082B94, 
                              32'h70486858, 32'h8F45FD19, 32'h94DE6C87, 32'h527BF8B7, 32'hAB73D323, 32'h724B02E2, 32'hE31F8F57, 32'h6655AB2A, 32'hB2EB2807, 32'h2FB5C203, 32'h86C57B9A, 32'hD33708A5, 32'h302887F2, 32'h23BFA5B2, 32'h02036ABA, 32'hED16825C, 
                              32'h8ACF1C2B, 32'hA779B492, 32'hF307F2F0, 32'h4E69E2A1, 32'h65DAF4CD, 32'h0605BED5, 32'hD134621F, 32'hC4A6FE8A, 32'h342E539D, 32'hA2F355A0, 32'h058AE132, 32'hA4F6EB75, 32'h0B83EC39, 32'h4060EFAA, 32'h5E719F06, 32'hBD6E1051, 
                              32'h3E218AF9, 32'h96DD063D, 32'hDD3E05AE, 32'h4DE6BD46, 32'h91548DB5, 32'h71C45D05, 32'h0406D46F, 32'h605015FF, 32'h1998FB24, 32'hD6BDE997, 32'h894043CC, 32'h67D99E77, 32'hB0E842BD, 32'h07898B88, 32'hE7195B38, 32'h79C8EEDB, 
                              32'hA17C0A47, 32'h7C420FE9, 32'hF8841EC9, 32'h00000000, 32'h09808683, 32'h322BED48, 32'h1E1170AC, 32'h6C5A724E, 32'hFD0EFFFB, 32'h0F853856, 32'h3DAED51E, 32'h362D3927, 32'h0A0FD964, 32'h685CA621, 32'h9B5B54D1, 32'h24362E3A, 
                              32'h0C0A67B1, 32'h9357E70F, 32'hB4EE96D2, 32'h1B9B919E, 32'h80C0C54F, 32'h61DC20A2, 32'h5A774B69, 32'h1C121A16, 32'hE293BA0A, 32'hC0A02AE5, 32'h3C22E043, 32'h121B171D, 32'h0E090D0B, 32'hF28BC7AD, 32'h2DB6A8B9, 32'h141EA9C8, 
                              32'h57F11985, 32'hAF75074C, 32'hEE99DDBB, 32'hA37F60FD, 32'hF701269F, 32'h5C72F5BC, 32'h44663BC5, 32'h5BFB7E34, 32'h8B432976, 32'hCB23C6DC, 32'hB6EDFC68, 32'hB8E4F163, 32'hD731DCCA, 32'h42638510, 32'h13972240, 32'h84C61120, 
                              32'h854A247D, 32'hD2BB3DF8, 32'hAEF93211, 32'hC729A16D, 32'h1D9E2F4B, 32'hDCB230F3, 32'h0D8652EC, 32'h77C1E3D0, 32'h2BB3166C, 32'hA970B999, 32'h119448FA, 32'h47E96422, 32'hA8FC8CC4, 32'hA0F03F1A, 32'h567D2CD8, 32'h223390EF, 
                              32'h87494EC7, 32'hD938D1C1, 32'h8CCAA2FE, 32'h98D40B36, 32'hA6F581CF, 32'hA57ADE28, 32'hDAB78E26, 32'h3FADBFA4, 32'h2C3A9DE4, 32'h5078920D, 32'h6A5FCC9B, 32'h547E4662, 32'hF68D13C2, 32'h90D8B8E8, 32'h2E39F75E, 32'h82C3AFF5, 
                              32'h9F5D80BE, 32'h69D0937C, 32'h6FD52DA9, 32'hCF2512B3, 32'hC8AC993B, 32'h10187DA7, 32'hE89C636E, 32'hDB3BBB7B, 32'hCD267809, 32'h6E5918F4, 32'hEC9AB701, 32'h834F9AA8, 32'hE6956E65, 32'hAAFFE67E, 32'h21BCCF08, 32'hEF15E8E6, 
                              32'hBAE79BD9, 32'h4A6F36CE, 32'hEA9F09D4, 32'h29B07CD6, 32'h31A4B2AF, 32'h2A3F2331, 32'hC6A59430, 32'h35A266C0, 32'h744EBC37, 32'hFC82CAA6, 32'hE090D0B0, 32'h33A7D815, 32'hF104984A, 32'h41ECDAF7, 32'h7FCD500E, 32'h1791F62F, 
                              32'h764DD68D, 32'h43EFB04D, 32'hCCAA4D54, 32'hE49604DF, 32'h9ED1B5E3, 32'h4C6A881B, 32'hC12C1FB8, 32'h4665517F, 32'h9D5EEA04, 32'h018C355D, 32'hFA877473, 32'hFB0B412E, 32'hB3671D5A, 32'h92DBD252, 32'hE9105633, 32'h6DD64713, 
                              32'h9AD7618C, 32'h37A10C7A, 32'h59F8148E, 32'hEB133C89, 32'hCEA927EE, 32'hB761C935, 32'hE11CE5ED, 32'h7A47B13C, 32'h9CD2DF59, 32'h55F2733F, 32'h1814CE79, 32'h73C737BF, 32'h53F7CDEA, 32'h5FFDAA5B, 32'hDF3D6F14, 32'h7844DB86, 
                              32'hCAAFF381, 32'hB968C43E, 32'h3824342C, 32'hC2A3405F, 32'h161DC372, 32'hBCE2250C, 32'h283C498B, 32'hFF0D9541, 32'h39A80171, 32'h080CB3DE, 32'hD8B4E49C, 32'h6456C190, 32'h7BCB8461, 32'hD532B670, 32'h486C5C74, 32'hD0B85742, 
                              // Inv_S_box
                                    // 0          1             2             3              4             5            6              7             8            9              A           B              C             D             E                                                                  
					32'h52000000, 32'h09000000, 32'h6a000000, 32'hd5000000, 32'h30000000, 32'h36000000, 32'ha5000000, 32'h38000000, 32'hbf000000, 32'h40000000, 32'ha3000000, 32'h9e000000, 32'h81000000, 32'hf3000000, 32'hd7000000, 32'hfb000000, 
                              32'h7c000000, 32'he3000000, 32'h39000000, 32'h82000000, 32'h9b000000, 32'h2f000000, 32'hff000000, 32'h87000000, 32'h34000000, 32'h8e000000, 32'h43000000, 32'h44000000, 32'hc4000000, 32'hde000000, 32'he9000000, 32'hcb000000, 
                              32'h54000000, 32'h7b000000, 32'h94000000, 32'h32000000, 32'ha6000000, 32'hc2000000, 32'h23000000, 32'h3d000000, 32'hee000000, 32'h4c000000, 32'h95000000, 32'h0b000000, 32'h42000000, 32'hfa000000, 32'hc3000000, 32'h4e000000, 
                              32'h08000000, 32'h2e000000, 32'ha1000000, 32'h66000000, 32'h28000000, 32'hd9000000, 32'h24000000, 32'hb2000000, 32'h76000000, 32'h5b000000, 32'ha2000000, 32'h49000000, 32'h6d000000, 32'h8b000000, 32'hd1000000, 32'h25000000, 
                              32'h72000000, 32'hf8000000, 32'hf6000000, 32'h64000000, 32'h86000000, 32'h68000000, 32'h98000000, 32'h16000000, 32'hd4000000, 32'ha4000000, 32'h5c000000, 32'hcc000000, 32'h5d000000, 32'h65000000, 32'hb6000000, 32'h92000000, 
                              32'h6c000000, 32'h70000000, 32'h48000000, 32'h50000000, 32'hfd000000, 32'hed000000, 32'hb9000000, 32'hda000000, 32'h5e000000, 32'h15000000, 32'h46000000, 32'h57000000, 32'ha7000000, 32'h8d000000, 32'h9d000000, 32'h84000000, 
                              32'h90000000, 32'hd8000000, 32'hab000000, 32'h00000000, 32'h8c000000, 32'hbc000000, 32'hd3000000, 32'h0a000000, 32'hf7000000, 32'he4000000, 32'h58000000, 32'h05000000, 32'hb8000000, 32'hb3000000, 32'h45000000, 32'h06000000, 
                              32'hd0000000, 32'h2c000000, 32'h1e000000, 32'h8f000000, 32'hca000000, 32'h3f000000, 32'h0f000000, 32'h02000000, 32'hc1000000, 32'haf000000, 32'hbd000000, 32'h03000000, 32'h01000000, 32'h13000000, 32'h8a000000, 32'h6b000000, 
                              32'h3a000000, 32'h91000000, 32'h11000000, 32'h41000000, 32'h4f000000, 32'h67000000, 32'hdc000000, 32'hea000000, 32'h97000000, 32'hf2000000, 32'hcf000000, 32'hce000000, 32'hf0000000, 32'hb4000000, 32'he6000000, 32'h73000000, 
                              32'h96000000, 32'hac000000, 32'h74000000, 32'h22000000, 32'he7000000, 32'had000000, 32'h35000000, 32'h85000000, 32'he2000000, 32'hf9000000, 32'h37000000, 32'he8000000, 32'h1c000000, 32'h75000000, 32'hdf000000, 32'h6e000000, 
                              32'h47000000, 32'hf1000000, 32'h1a000000, 32'h71000000, 32'h1d000000, 32'h29000000, 32'hc5000000, 32'h89000000, 32'h6f000000, 32'hb7000000, 32'h62000000, 32'h0e000000, 32'haa000000, 32'h18000000, 32'hbe000000, 32'h1b000000, 
                              32'hfc000000, 32'h56000000, 32'h3e000000, 32'h4b000000, 32'hc6000000, 32'hd2000000, 32'h79000000, 32'h20000000, 32'h9a000000, 32'hdb000000, 32'hc0000000, 32'hfe000000, 32'h78000000, 32'hcd000000, 32'h5a000000, 32'hf4000000, 
                              32'h1f000000, 32'hdd000000, 32'ha8000000, 32'h33000000, 32'h88000000, 32'h07000000, 32'hc7000000, 32'h31000000, 32'hb1000000, 32'h12000000, 32'h10000000, 32'h59000000, 32'h27000000, 32'h80000000, 32'hec000000, 32'h5f000000, 
                              32'h60000000, 32'h51000000, 32'h7f000000, 32'ha9000000, 32'h19000000, 32'hb5000000, 32'h4a000000, 32'h0d000000, 32'h2d000000, 32'he5000000, 32'h7a000000, 32'h9f000000, 32'h93000000, 32'hc9000000, 32'h9c000000, 32'hef000000, 
                              32'ha0000000, 32'he0000000, 32'h3b000000, 32'h4d000000, 32'hae000000, 32'h2a000000, 32'hf5000000, 32'hb0000000, 32'hc8000000, 32'heb000000, 32'hbb000000, 32'h3c000000, 32'h83000000, 32'h53000000, 32'h99000000, 32'h61000000, 
                              32'h17000000, 32'h2b000000, 32'h04000000, 32'h7e000000, 32'hba000000, 32'h77000000, 32'hd6000000, 32'h26000000, 32'he1000000, 32'h69000000, 32'h14000000, 32'h63000000, 32'h55000000, 32'h21000000, 32'h0c000000, 32'h7d000000
                              };
									
always_comb begin
      if(!i_reset) begin
            o_data = 32'h0;
      end
      else
      begin
            o_data = mem[address];
      end
end		 

endmodule 

`endif